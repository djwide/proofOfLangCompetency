-------------------------------------------------------------------------------
-- EE375 Datapath for MARC2 Processor
-- Author:         David Weidman
-- Date Modified:  26 JAN 15
-------------------------------------------------------------------------------


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY datapath IS
  PORT( clk: IN std_logic; 	    -- clock	
        rst : IN STD_LOGIC;		
        rWE: IN std_logic;      -- register file & flag write enable
        ld_op: IN std_logic;	-- op is load (from control unit)
        st_op: IN std_logic; 	-- op is store (from control unit)
        ctlWd: IN  std_logic_vector(14 downto 0);    -- control word
        const_in: IN  std_logic_vector(15 downto 0); -- data from control unit
        N: OUT std_logic; 	-- negative flag (N=1, sign of result is neg)
        Z: OUT std_logic; 	-- zero flag (Z=1, result of Func Unit is 0)
        R0out,R1out,R2out,R3out, R4out,R5out,R6out,R7out: OUT std_logic_vector(15 downto 0);
        dp_addr_bus: OUT std_logic_vector(15 downto 0);    -- address to memory
        dp_data_bus: INOUT std_logic_vector(15 downto 0)); -- data to/from memory
END datapath;

ARCHITECTURE DPArch OF datapath IS
------------------------------------------------------------------------------- 
-- control word format
--      |cw(14)|cw(13)|cw(12-10)|cw(9-6)|cw(5-3)|cw(2-0)| 
--      |  MD  |  MB  |  selD   |  FS   |  selA |  selB |
-------------------------------------------------------------------------------
  -- component declarations
		
	component regFile is
		PORT( clk: IN std_logic; 	    
		  rst : IN STD_LOGIC;		
		  rWE: IN std_logic;    
		  dataIn: IN  std_logic_vector(15 downto 0);    
		  ctlWd: IN  std_logic_vector(14 downto 0);  
		  R0out,R1out,R2out,R3out,R4out,R5out,R6out,R7out: OUT std_logic_vector(15 downto 0);
		  A_bus: OUT std_logic_vector(15 downto 0);   
		  B_bus: INOUT std_logic_vector(15 downto 0)); 
		  --Hwang, Colin CDT H-2 '16.  Assistance given to author verbally confirming that a semicolon is 
		  --not in fact needed between the parentheses as well as after the parentheses.
		  -- This same piece of syntax applies to the port declarations in the components as well
		end component;
		
	component mux2_1 is
		PORT(a,b: IN std_logic_vector(15 downto 0);
			s: IN std_logic;
			y: out std_logic_vector(15 downto 0));
	end component;
	
	Component ALU is
		PORT(A,B: IN std_logic_vector(15 downto 0);
			sel: IN std_logic_vector(3 downto 0);
			F: buffer std_logic_vector(15 downto 0);
			Z, N: OUT std_logic);
		end component;
	
	component triStateBuffer is 
		port(A: in Std_logic_vector(15 downto 0);
		A_En: in STD_Logic;
		F: out Std_logic_vector(15 downto 0));
	end component;
			
	signal aInput: std_logic;
	SIGNAL aBus, bBus,bRFOut,aluOut,rfIn : std_logic_vector(15 DOWNTO 0);
  
BEGIN 
	regF: regFile PORT MAP(clk,rst,rWE,rfIn,ctlWd,R0out,R1out,R2out,R3out,R4out,R5out,R6out,R7out,aBus,bRFOut);
	ALU1 : ALU PORT MAP(aBus,bBus,ctlWd(9 downto 6), aluOut, Z, N);
	MD : mux2_1 PORT MAP(aluOut,dp_data_bus,ctlWd(14), rfIn);
	MB : mux2_1 PORT MAP(bRFOut,const_in,ctlWd(13), bBus);
	TSBA : triStateBuffer PORT MAP(aBus,aInput,dp_addr_bus);
	TSBB : triStateBuffer PORT MAP(bBus,st_op,dp_data_bus);
	aInput <= ld_op or st_op;
END DPArch;