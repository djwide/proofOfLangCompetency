--------------------------------------------------------------------------------------		
--	File:  CPU_chip.vhd
--	Created by: MAJ Paul Maxwell
--	Date Created:  4 Sep 03
--	Modified by:  MAJ Julianna Rodriguez
--	Date Last Modified:  20150217
-- 	Description:  This file provides the top-level design for the EE375 MARC2 
--			processor.  Using the constraints file provided and this code, the user can
--			insert a cadet's MARC2 source code into this project (replacing my cpu_marc1
--			and its dependent files) and implement this processor in hardware.  This 
--			solution is designed for an Altera Cyclone IVE chip on an 
--			Terasic DE2-115 Education and Development Board.  
-------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CPU_chip is
    Port( clk : in std_logic;                              -- CPU clock
          reset : in std_logic;                            -- key0
          run : in std_logic;                              -- SW17 
          reg_select : in STD_LOGIC_VECTOR(2 downto 0);    -- SW2-SW0 select lines for register output
          LCD_RS, LCD_E, LCD_ON: out std_logic;   				-- lcd control signals
          LCD_RW   :buffer std_logic;
			 rstLED, prgmLED : out std_logic;                 -- led drivers
          lcd_data : INOUT	STD_LOGIC_VECTOR(7 DOWNTO 0)); -- data lines to lcd displayReg
end CPU_chip;



architecture Behavioral of CPU_chip is
  COMPONENT CPU IS
    PORT( clk, reset, run           : IN std_logic;				
          mem_rd, mem_wr          : OUT std_logic;	
          address             	 : OUT std_logic_vector(15 downto 0);
          R0out,R1out,R2out,R3out : OUT std_logic_vector(15 downto 0);  
          R4out,R5out,R6out,R7out : OUT std_logic_vector(15 downto 0);
			 data							 : INOUT std_logic_vector(15 downto 0));
  END COMPONENT;

-- The following RAM and ROM are generated by the Coregen tool.  They are created as
-- single port block memory units which are clocked on the falling edge in order to 
-- remove some timing conflicts.
  COMPONENT systemROM IS
	PORT( address : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		   clock	  : IN STD_LOGIC  := '1';
		   q       : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
  END COMPONENT;

  COMPONENT systemRAM IS
	PORT( address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
		   clock	  : IN STD_LOGIC  := '1';
		   data    : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		   wren    : IN STD_LOGIC ;
		   q       : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
  END COMPONENT;

  COMPONENT LCDdisplay IS
    PORT( reset, clk_50Mhz              : IN STD_LOGIC;
          LCD_RS, LCD_E, LCD_ON, rstLED : OUT STD_LOGIC;
          LCD_RW                        : BUFFER STD_LOGIC;
          display_data                  : IN STD_LOGIC_VECTOR(15 downto 0);
          DATA_BUS                      : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0));
  END COMPONENT;
  
signal mem_rd, mem_wr, lcdRW : std_logic;
signal Addr_bus, Data_bus, ROM_data, RAM_data : std_logic_vector(15 downto 0);
signal R0out,R1out,R2out,R3out,R4out,R5out,R6out,R7out : std_logic_vector(15 downto 0);
signal DisplayReg, display_buf : std_logic_vector(15 downto 0);

begin
prgmLED <= '1';

Data_bus <= ROM_data when (mem_rd='1' and addr_bus(15 downto 12)="0000") else
            RAM_data when (mem_rd='1') else
            (others=>'Z');	  

displayReg <= R0out when reg_select = "000" else
              R1out when reg_select = "001" else
              R2out when reg_select = "010" else
              R3out when reg_select = "011" else
              R4out when reg_select = "100" else
              R5out when reg_select = "101" else	
              R6out when reg_select = "110" else
              R7out when reg_select = "111" else
              x"F0BA";    -- short for FUBAR                  
				  
RAM1 : systemRAM port map (address=>addr_bus(14 downto 0), clock=>clk, 
                           data=>Data_bus, wren=>mem_wr, q=>RAM_data);

ROM1 : systemROM port map (address=>addr_bus(11 downto 0), clock=>clk, 
                           q=>ROM_data);

CPU1: CPU port map(clk=>clk, reset=>reset, run=>run,
						mem_rd=>mem_rd, mem_wr=>mem_wr, address=>addr_bus, 
                   R0out=>R0out, R1out=>R1out, R2out=>R2out, R3out=>R3out,
                   R4out=>R4out, R5out=>R5out, R6out=>R6out, R7out=>R7out,
						 data=>Data_bus); 	
			
lcd_out: LCDdisplay port map( reset, clk, LCD_RS, LCD_E, LCD_ON, rstLED, LCD_RW, 
                              displayReg, lcd_data);
		  
end Behavioral;
